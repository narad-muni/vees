module main

struct Driver{

}

struct ChromeDriver{

}

struct Element{
	
}

fn main() {
	println('Hello World!')
}
